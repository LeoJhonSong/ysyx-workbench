// 双控开关, ysyx预学习0.4
module top(
  input a,
  input b,
  output f
);
  assign f = a ^ b;
endmodule
